 module mips_tb();
    
   reg clk, rst;
    
   mips U_MIPS(
      .clk(clk), .rst(rst)
   );
    
    initial begin
        // $readmemh("Test_6_Instr.txt" , U_MIPS.U_IM.imem) ;
        $readmemh("test.txt" , U_MIPS.U_IM.imem) ;
        $monitor("        PC = 0x%8X\n        IR = 0x%8X", U_MIPS.U_PC.PC, U_MIPS.U_IM.dout);
        
        clk = 1 ;
        rst = 0 ;
        #5 ;
        rst = 1 ;
        #20 ;
        rst = 0 ;
    end

    always
    #(50) clk = ~clk;
endmodule
